//Copyright (C)2014-2024 Gowin Semiconductor Corporation.
//All rights reserved.
//File Title: IP file
//Tool Version: V1.9.9.02
//Part Number: GW1NZ-LV1QN48A3
//Device: GW1NZ-1
//Device Version: C
//Created Time: Wed Jul 17 21:54:29 2024

module charBuffer (dout, clk, oce, ce, reset, wre, ad, din);

output [7:0] dout;
input clk;
input oce;
input ce;
input reset;
input wre;
input [11:0] ad;
input [7:0] din;

wire [27:0] sp_inst_0_dout_w;
wire [27:0] sp_inst_1_dout_w;
wire gw_gnd;

assign gw_gnd = 1'b0;

SP sp_inst_0 (
    .DO({sp_inst_0_dout_w[27:0],dout[3:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,gw_gnd}),
    .AD({ad[11:0],gw_gnd,gw_gnd}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[3:0]})
);

defparam sp_inst_0.READ_MODE = 1'b0;
defparam sp_inst_0.WRITE_MODE = 2'b10;
defparam sp_inst_0.BIT_WIDTH = 4;
defparam sp_inst_0.BLK_SEL = 3'b000;
defparam sp_inst_0.RESET_MODE = "SYNC";
defparam sp_inst_0.INIT_RAM_00 = 256'h0;
defparam sp_inst_0.INIT_RAM_01 = 256'h0;
defparam sp_inst_0.INIT_RAM_02 = 256'h0;
defparam sp_inst_0.INIT_RAM_03 = 256'h0;
defparam sp_inst_0.INIT_RAM_04 = 256'h0;
defparam sp_inst_0.INIT_RAM_05 = 256'h0;
defparam sp_inst_0.INIT_RAM_06 = 256'h0;
defparam sp_inst_0.INIT_RAM_07 = 256'h0;
defparam sp_inst_0.INIT_RAM_08 = 256'h0;
defparam sp_inst_0.INIT_RAM_09 = 256'h0;
defparam sp_inst_0.INIT_RAM_0A = 256'h0;
defparam sp_inst_0.INIT_RAM_0B = 256'h0;
defparam sp_inst_0.INIT_RAM_0C = 256'h0;
defparam sp_inst_0.INIT_RAM_0D = 256'h0;
defparam sp_inst_0.INIT_RAM_0E = 256'h0;
defparam sp_inst_0.INIT_RAM_0F = 256'h0;
defparam sp_inst_0.INIT_RAM_10 = 256'h0;
defparam sp_inst_0.INIT_RAM_11 = 256'h0;
defparam sp_inst_0.INIT_RAM_12 = 256'h0;
defparam sp_inst_0.INIT_RAM_13 = 256'h0;
defparam sp_inst_0.INIT_RAM_14 = 256'h0;
defparam sp_inst_0.INIT_RAM_15 = 256'h0;
defparam sp_inst_0.INIT_RAM_16 = 256'h0;
defparam sp_inst_0.INIT_RAM_17 = 256'h0;
defparam sp_inst_0.INIT_RAM_18 = 256'h0;
defparam sp_inst_0.INIT_RAM_19 = 256'h0;
defparam sp_inst_0.INIT_RAM_1A = 256'h0;
defparam sp_inst_0.INIT_RAM_1B = 256'h0;
defparam sp_inst_0.INIT_RAM_1C = 256'h0;
defparam sp_inst_0.INIT_RAM_1D = 256'h0;
defparam sp_inst_0.INIT_RAM_1E = 256'h0;
defparam sp_inst_0.INIT_RAM_1F = 256'h0;
defparam sp_inst_0.INIT_RAM_20 = 256'h0;
defparam sp_inst_0.INIT_RAM_21 = 256'h0;
defparam sp_inst_0.INIT_RAM_22 = 256'h0;
defparam sp_inst_0.INIT_RAM_23 = 256'h0;
defparam sp_inst_0.INIT_RAM_24 = 256'h0;
defparam sp_inst_0.INIT_RAM_25 = 256'h0;
defparam sp_inst_0.INIT_RAM_26 = 256'h0;
defparam sp_inst_0.INIT_RAM_27 = 256'h0;

SP sp_inst_1 (
    .DO({sp_inst_1_dout_w[27:0],dout[7:4]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,gw_gnd}),
    .AD({ad[11:0],gw_gnd,gw_gnd}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[7:4]})
);

defparam sp_inst_1.READ_MODE = 1'b0;
defparam sp_inst_1.WRITE_MODE = 2'b10;
defparam sp_inst_1.BIT_WIDTH = 4;
defparam sp_inst_1.BLK_SEL = 3'b000;
defparam sp_inst_1.RESET_MODE = "SYNC";
defparam sp_inst_1.INIT_RAM_00 = 256'h0;
defparam sp_inst_1.INIT_RAM_01 = 256'h0;
defparam sp_inst_1.INIT_RAM_02 = 256'h0;
defparam sp_inst_1.INIT_RAM_03 = 256'h0;
defparam sp_inst_1.INIT_RAM_04 = 256'h0;
defparam sp_inst_1.INIT_RAM_05 = 256'h0;
defparam sp_inst_1.INIT_RAM_06 = 256'h0;
defparam sp_inst_1.INIT_RAM_07 = 256'h0;
defparam sp_inst_1.INIT_RAM_08 = 256'h0;
defparam sp_inst_1.INIT_RAM_09 = 256'h0;
defparam sp_inst_1.INIT_RAM_0A = 256'h0;
defparam sp_inst_1.INIT_RAM_0B = 256'h0;
defparam sp_inst_1.INIT_RAM_0C = 256'h0;
defparam sp_inst_1.INIT_RAM_0D = 256'h0;
defparam sp_inst_1.INIT_RAM_0E = 256'h0;
defparam sp_inst_1.INIT_RAM_0F = 256'h0;
defparam sp_inst_1.INIT_RAM_10 = 256'h0;
defparam sp_inst_1.INIT_RAM_11 = 256'h0;
defparam sp_inst_1.INIT_RAM_12 = 256'h0;
defparam sp_inst_1.INIT_RAM_13 = 256'h0;
defparam sp_inst_1.INIT_RAM_14 = 256'h0;
defparam sp_inst_1.INIT_RAM_15 = 256'h0;
defparam sp_inst_1.INIT_RAM_16 = 256'h0;
defparam sp_inst_1.INIT_RAM_17 = 256'h0;
defparam sp_inst_1.INIT_RAM_18 = 256'h0;
defparam sp_inst_1.INIT_RAM_19 = 256'h0;
defparam sp_inst_1.INIT_RAM_1A = 256'h0;
defparam sp_inst_1.INIT_RAM_1B = 256'h0;
defparam sp_inst_1.INIT_RAM_1C = 256'h0;
defparam sp_inst_1.INIT_RAM_1D = 256'h0;
defparam sp_inst_1.INIT_RAM_1E = 256'h0;
defparam sp_inst_1.INIT_RAM_1F = 256'h0;
defparam sp_inst_1.INIT_RAM_20 = 256'h0;
defparam sp_inst_1.INIT_RAM_21 = 256'h0;
defparam sp_inst_1.INIT_RAM_22 = 256'h0;
defparam sp_inst_1.INIT_RAM_23 = 256'h0;
defparam sp_inst_1.INIT_RAM_24 = 256'h0;
defparam sp_inst_1.INIT_RAM_25 = 256'h0;
defparam sp_inst_1.INIT_RAM_26 = 256'h0;
defparam sp_inst_1.INIT_RAM_27 = 256'h0;

endmodule //charBuffer
