//Copyright (C)2014-2024 Gowin Semiconductor Corporation.
//All rights reserved.
//File Title: IP file
//Tool Version: V1.9.9.02
//Part Number: GW1NZ-LV1QN48C6/I5
//Device: GW1NZ-1
//Created Time: Sun Jun 15 21:30:12 2025

module charROM (dout, clk, oce, ce, reset, ad);

output [7:0] dout;
input clk;
input oce;
input ce;
input reset;
input [10:0] ad;

wire [23:0] prom_inst_0_dout_w;
wire gw_gnd;

assign gw_gnd = 1'b0;

pROM prom_inst_0 (
    .DO({prom_inst_0_dout_w[23:0],dout[7:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .AD({ad[10:0],gw_gnd,gw_gnd,gw_gnd})
);

defparam prom_inst_0.READ_MODE = 1'b0;
defparam prom_inst_0.BIT_WIDTH = 8;
defparam prom_inst_0.RESET_MODE = "SYNC";
defparam prom_inst_0.INIT_RAM_00 = 256'h007E080800000E0000880008000000A000000400A00000000C81160018A89000;
defparam prom_inst_0.INIT_RAM_01 = 256'h3E10000400001E1E3F1E3F021E1E081E00000000000008081018200812120800;
defparam prom_inst_0.INIT_RAM_02 = 256'h00081C001C3F21212122217F1E3E1C3E0C214120211F3E211E3F3F3E1E3E0C3E;
defparam prom_inst_0.INIT_RAM_03 = 256'h3E3038100E00A10000000000000082A00000001040B80040C20C000200400002;
defparam prom_inst_0.INIT_RAM_04 = 256'h3020081C0000101C00880008000000A000000E00A070000012810E0024A89000;
defparam prom_inst_0.INIT_RAM_05 = 256'h4108000800002121212120062121182101000000080004101014503E12120800;
defparam prom_inst_0.INIT_RAM_06 = 256'h0014044010012121212221082121222112316320220408212120201121111241;
defparam prom_inst_0.INIT_RAM_07 = 256'h3E49041010009E0000000010000083A00000001040040840BC12000200400002;
defparam prom_inst_0.INIT_RAM_08 = 256'h4910082A100410220000003E0000000040001000001820002100101820900000;
defparam prom_inst_0.INIT_RAM_09 = 256'h61040010181821210220200A0101282102000000084902202014224812120800;
defparam prom_inst_0.INIT_RAM_0A = 256'h002204201002211221222108202122212129552024040821402020112011214D;
defparam prom_inst_0.INIT_RAM_0B = 256'h3E06041010000000000000100000000000000010400000400010000200400001;
defparam prom_inst_0.INIT_RAM_0C = 256'h060808082002102222490149323F1F1E3F0C0C31241C24102116202010610E00;
defparam prom_inst_0.INIT_RAM_0D = 256'h02023F2000002121042020120102082304000000082A0220001404487F000800;
defparam prom_inst_0.INIT_RAM_0E = 256'h004104101004120C212221082021222121294920280408214020201120112153;
defparam prom_inst_0.INIT_RAM_0F = 256'h3E000400103F21214122427C3C2E1E3E3C2E7610440418583E103C3A3C5C3C00;
defparam prom_inst_0.INIT_RAM_10 = 256'h000408087F7F1022414962491248242112121011241228103F2940401C121119;
defparam prom_inst_0.INIT_RAM_11 = 256'h0C01004000001F1E083E3E220E04082508003F007F1C02200008083E12000800;
defparam prom_inst_0.INIT_RAM_12 = 256'h0000040810080C0C212221081E3E223E212549203004083F403C3C11201E3F51;
defparam prom_inst_0.INIT_RAM_13 = 256'h3E0002002002211249224210423122214231491048040864427C424642620200;
defparam prom_inst_0.INIT_RAM_14 = 256'h3008080820021022494914491208422112212012241230102109407824141F25;
defparam prom_inst_0.INIT_RAM_15 = 256'h10023F20180001210821013F0108082910000018081C0220001510097F000800;
defparam prom_inst_0.INIT_RAM_16 = 256'h000004041010040C2D2221080128222021234120280408214720201120112152;
defparam prom_inst_0.INIT_RAM_17 = 256'h3E0004101004210C492242103020222142214910700408424210424240423E00;
defparam prom_inst_0.INIT_RAM_18 = 256'h49102A0810045014494A083E1208422212211E14241228102109384024181122;
defparam prom_inst_0.INIT_RAM_19 = 256'h1004001008180121082101020110083120000008082A02200022240912000000;
defparam prom_inst_0.INIT_RAM_1A = 256'h00000402102004122D22210801242A202123412024040821412020112011214C;
defparam prom_inst_0.INIT_RAM_1B = 256'h3E0004101008230C492242100C202231422149104804084246107E4240424200;
defparam prom_inst_0.INIT_RAM_1C = 256'h06201C0800003014493C14081208243C121201183A1225141209042024101E25;
defparam prom_inst_0.INIT_RAM_1D = 256'h00080008080021210821210221200821401800080849041000224A7E12000000;
defparam prom_inst_0.INIT_RAM_1E = 256'h0000040110200421331421082122262012214120224408212120201121112141;
defparam prom_inst_0.INIT_RAM_1F = 256'h3E00041010101D124914421242203E2E42214910440408423A10404642624600;
defparam prom_inst_0.INIT_RAM_20 = 256'h007E080800001036360823080E081820130C06102033220C0C01181818281019;
defparam prom_inst_0.INIT_RAM_21 = 256'h1810000410001E1E081E1E021E3F3E1E0018001000000808001D040812000800;
defparam prom_inst_0.INIT_RAM_22 = 256'h7F001C001C3F042121081E081E211D200C21413E21383E211E203F3E1E3E213E;
defparam prom_inst_0.INIT_RAM_23 = 256'h3E0038000E3F012136083C0C3C2002203C21490C42440C4202103E3A3C5C3B00;

endmodule //charROM
