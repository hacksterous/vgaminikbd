	`ifdef SIM_ONLY
	`define DELAY #1
	`else
	`define DELAY 
	`endif
	//`define DEBUG_FPGA_BUILD
	`undef DEBUG_FPGA_BUILD
