//Copyright (C)2014-2024 Gowin Semiconductor Corporation.
//All rights reserved.
//File Title: IP file
//Tool Version: V1.9.9.02
//Part Number: GW1NZ-LV1QN48A3
//Device: GW1NZ-1
//Device Version: C
//Created Time: Wed Jul 17 20:29:19 2024

module charROM (dout, clk, oce, ce, reset, ad);

output [4:0] dout;
input clk;
input oce;
input ce;
input reset;
input [10:0] ad;

wire [26:0] prom_inst_0_dout_w;
wire gw_gnd;

assign gw_gnd = 1'b0;

pROM prom_inst_0 (
    .DO({prom_inst_0_dout_w[26:0],dout[4:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .AD({ad[10:0],gw_gnd,gw_gnd,gw_gnd})
);

defparam prom_inst_0.READ_MODE = 1'b0;
defparam prom_inst_0.BIT_WIDTH = 8;
defparam prom_inst_0.RESET_MODE = "SYNC";
defparam prom_inst_0.INIT_RAM_00 = 256'h00040E1F1F1F0A00000E1B111F151F0E000E111B1F151F0E0000000000000000;
defparam prom_inst_0.INIT_RAM_01 = 256'h0000040E0E040000000E041F1F1F0E04000E041F151F0A0E00040E1F1F0E0400;
defparam prom_inst_0.INIT_RAM_02 = 256'h000814140D0307001F1F1B15151B1F1F0000040A0A0400001F1F1B11111B1F1F;
defparam prom_inst_0.INIT_RAM_03 = 256'h04150E1B1B0E150400180B09090F090F00180808080F090F00041F040E11110E;
defparam prom_inst_0.INIT_RAM_04 = 256'h001B001B1B1B1B1B00040E1504150E040001030F1F0F03010010181E1F1E1810;
defparam prom_inst_0.INIT_RAM_05 = 256'h1F040E1504150E04001F1F000000000006090902050A0906000505050D15150F;
defparam prom_inst_0.INIT_RAM_06 = 256'h000004081F080400000004021F02040000040E150404040000040404150E0400;
defparam prom_inst_0.INIT_RAM_07 = 256'h000004040E1F1F0000001F1F0E0404000000000A1F1F0A000000001F10101000;
defparam prom_inst_0.INIT_RAM_08 = 256'h000A0A1F0A1F0A0A00000000000A0A0A00040004040404040000000000000000;
defparam prom_inst_0.INIT_RAM_09 = 256'h0000000008040606000D121508141408000313080402191800041E050E140F04;
defparam prom_inst_0.INIT_RAM_0A = 256'h000004041F0404000004150E1F0E150400080402020204080002040808080402;
defparam prom_inst_0.INIT_RAM_0B = 256'h00001008040201000006060000000000000000001F0000000804060600000000;
defparam prom_inst_0.INIT_RAM_0C = 256'h000E11010602011F001F10100E01110E000E040404040C04000E11191513110E;
defparam prom_inst_0.INIT_RAM_0D = 256'h001008040201011F000E11111E100807000E1101011E101F0002021F120A0602;
defparam prom_inst_0.INIT_RAM_0E = 256'h00080404000400000000000400040000001C02010F11110E000E11110E11110E;
defparam prom_inst_0.INIT_RAM_0F = 256'h000400040601110E00080402010204080000001F001F00000001020408040201;
defparam prom_inst_0.INIT_RAM_10 = 256'h000E11101010110E001E11111E11111E0011111F11110A04000F10161715110E;
defparam prom_inst_0.INIT_RAM_11 = 256'h000F11131010110F001010101E10101F001F10101E10101F001E11111111111E;
defparam prom_inst_0.INIT_RAM_12 = 256'h0011121418141211000C120202020207000E04040404040E001111111F111111;
defparam prom_inst_0.INIT_RAM_13 = 256'h000E11111111110E00111113151911110011111515151B11001F101010101010;
defparam prom_inst_0.INIT_RAM_14 = 256'h000E11010E10110E001112141E11111E000D12151111110E001010101E11111E;
defparam prom_inst_0.INIT_RAM_15 = 256'h000A15151511111100040A1111111111000E111111111111000404040404151F;
defparam prom_inst_0.INIT_RAM_16 = 256'h000F08080808080F001F10080E02011F00040404040A11110011110A040A1111;
defparam prom_inst_0.INIT_RAM_17 = 256'h001F0000000000000000000000110A04000F01010101010F0000010204081000;
defparam prom_inst_0.INIT_RAM_18 = 256'h000E1110110E00000016191119161010000F120E020C00000000000002040C0C;
defparam prom_inst_0.INIT_RAM_19 = 256'h0E010D13130E0000000404040E040502000E101F110E0000000D1311130D0101;
defparam prom_inst_0.INIT_RAM_1A = 256'h0012141814121010000C120202020002000E0404040C00040011111119161010;
defparam prom_inst_0.INIT_RAM_1B = 256'h000E1111110E0000001111111916000000151515151A0000000E04040404040C;
defparam prom_inst_0.INIT_RAM_1C = 256'h001E010E100F0000001010101916000001010D13130D00001010161919160000;
defparam prom_inst_0.INIT_RAM_1D = 256'h000A15151111000000040A1111110000000D13111111000000020504041F0404;
defparam prom_inst_0.INIT_RAM_1E = 256'h0002040408040402001F0804021F00000E11010F1111000000110A040A110000;
defparam prom_inst_0.INIT_RAM_1F = 256'h00001F11111B0E04000000000002150800080404020404080004040400040404;
defparam prom_inst_0.INIT_RAM_20 = 256'h000F120E020C001F000F101F110E0003000D1311110011000C020E111010110E;
defparam prom_inst_0.INIT_RAM_21 = 256'h0006020F18180F00000F120E020C0006000F120E020C0018000F120E020C0011;
defparam prom_inst_0.INIT_RAM_22 = 256'h0007020202060005000F101F110E0018000F101F110E0011000F101F110E001F;
defparam prom_inst_0.INIT_RAM_23 = 256'h11111F110A04000411111F110A04000A000702020206000C0007020202060906;
defparam prom_inst_0.INIT_RAM_24 = 256'h000E11110E00110E001312121F120A07000F120F020F0000001E101C101E0006;
defparam prom_inst_0.INIT_RAM_25 = 256'h000D131111001800000D13111100110E000E11110E001800000E11110E001100;
defparam prom_inst_0.INIT_RAM_26 = 256'h04041F14141F0404000E111111110011000E1111110E00110E01070909090009;
defparam prom_inst_0.INIT_RAM_27 = 256'h181404040E040503121217121C12121C04041F041F0E1B1B001F09081C090B06;
defparam prom_inst_0.INIT_RAM_28 = 256'h000D131111000300000E11110E0003000007020202060003000F120E020C0003;
defparam prom_inst_0.INIT_RAM_29 = 256'h00001F000E11110E00001F000F12120E001113171D19001F000909090E000F00;
defparam prom_inst_0.INIT_RAM_2A = 256'h0704130917121110000001011F000000000010101F000000000E11100C040004;
defparam prom_inst_0.INIT_RAM_2B = 256'h0000140A050A14000000050A140A050000040404040004040101170B15121110;
defparam prom_inst_0.INIT_RAM_2C = 256'h0202021E020202020202020202020202150A150A150A150A1104110411041104;
defparam prom_inst_0.INIT_RAM_2D = 256'h0202021E021E00000505051F000000000505051D050505050202021E021E0202;
defparam prom_inst_0.INIT_RAM_2E = 256'h0000001F011D05050505051D011F000005050505050505050505051D011D0505;
defparam prom_inst_0.INIT_RAM_2F = 256'h00000003020202020202021E000000000000001E021E02020000001F05050505;
defparam prom_inst_0.INIT_RAM_30 = 256'h0000001F0000000002020203020202020202021F000000000000001F02020202;
defparam prom_inst_0.INIT_RAM_31 = 256'h0000000704050505050505050505050502020203020302020202021F02020202;
defparam prom_inst_0.INIT_RAM_32 = 256'h05050505040505050505051D001F00000000001F001D05050505050504070000;
defparam prom_inst_0.INIT_RAM_33 = 256'h0000001F050505050000001F001F02020505051D001D05050000001F001F0000;
defparam prom_inst_0.INIT_RAM_34 = 256'h000000030203020200000007050505050505051F000000000202021F001F0000;
defparam prom_inst_0.INIT_RAM_35 = 256'h0202021F021F02020505051F0505050505050507000000000202020302030000;
defparam prom_inst_0.INIT_RAM_36 = 256'h1F1F1F1F000000001F1F1F1F1F1F1F1F02020203000000000000001E02020202;
defparam prom_inst_0.INIT_RAM_37 = 256'h000D1212120D0000000000001F1F1F1F03030303030303031C1C1C1C1C1C1C1C;
defparam prom_inst_0.INIT_RAM_38 = 256'h001F11080408111F000A0A0A0A0A1F000010101010131F0000101E131E130E00;
defparam prom_inst_0.INIT_RAM_39 = 256'h1F040E11110E041F0004040404141F0000180D0A0A0A0A00000C1212120F0000;
defparam prom_inst_0.INIT_RAM_3A = 256'h000E15150E000000000E11110E060806001B0A0A11110A0400040A111F110A04;
defparam prom_inst_0.INIT_RAM_3B = 256'h00001F001F001F00001111111111110E000E10101E10100E100E191515130E01;
defparam prom_inst_0.INIT_RAM_3C = 256'h0404040404040507001F000204080402001F000804020408001F0004041F0404;
defparam prom_inst_0.INIT_RAM_3D = 256'h000000000E1B1B0E0000171D00171D00000606001F0006061C14140404040404;
defparam prom_inst_0.INIT_RAM_3E = 256'h000000090909090E040C14140404040700000006000000000000000606000000;
defparam prom_inst_0.INIT_RAM_3F = 256'h0000000000000000000000000000000000000F0F0F0F00000000000F0C06030E;

endmodule //charROM
