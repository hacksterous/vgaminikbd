//Copyright (C)2014-2024 Gowin Semiconductor Corporation.
//All rights reserved.
//File Title: IP file
//Tool Version: V1.9.9.02
//Part Number: GW1NZ-LV1QN48C6/I5
//Device: GW1NZ-1
//Created Time: Fri May 30 18:41:38 2025

module charROM (dout, clk, oce, ce, reset, ad);

output [7:0] dout;
input clk;
input oce;
input ce;
input reset;
input [10:0] ad;

wire [23:0] prom_inst_0_dout_w;
wire gw_gnd;

assign gw_gnd = 1'b0;

pROM prom_inst_0 (
    .DO({prom_inst_0_dout_w[23:0],dout[7:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .AD({ad[10:0],gw_gnd,gw_gnd,gw_gnd})
);

defparam prom_inst_0.READ_MODE = 1'b0;
defparam prom_inst_0.BIT_WIDTH = 8;
defparam prom_inst_0.RESET_MODE = "SYNC";
defparam prom_inst_0.INIT_RAM_00 = 256'h007E080800000E0000880008000000A000000400A00000000C81160018909000;
defparam prom_inst_0.INIT_RAM_01 = 256'h3E10000400001E1E3F1E3F021E1E081E00000000000808081018200812120800;
defparam prom_inst_0.INIT_RAM_02 = 256'h00081C001C3F21212122217F1E3E1C3E0C214120211F3E211E3F3F3E1E3E0C3E;
defparam prom_inst_0.INIT_RAM_03 = 256'h3E3038100E00810000000000000082A00000001040840040820C000200400002;
defparam prom_inst_0.INIT_RAM_04 = 256'h3020081C0000101C00880008000000A000000E00A070000012810E0024909000;
defparam prom_inst_0.INIT_RAM_05 = 256'h41080008000021212121200621211821000000000C4904101014503E12120800;
defparam prom_inst_0.INIT_RAM_06 = 256'h0014044010012121212221082121222112316320220408212120201121111241;
defparam prom_inst_0.INIT_RAM_07 = 256'h3E4904101000A10000000010000082A00000001040C40840C212000200400002;
defparam prom_inst_0.INIT_RAM_08 = 256'h4910082A100410220088003E000000A040001000A01820002181101820909000;
defparam prom_inst_0.INIT_RAM_09 = 256'h61040010303021210220200A0101282101000000002A02202014224812120800;
defparam prom_inst_0.INIT_RAM_0A = 256'h002204201002211221222108202122212129552024040821402020112011215D;
defparam prom_inst_0.INIT_RAM_0B = 256'h3E06041010009E0000000010000083A00000001040B80040BC10000200400001;
defparam prom_inst_0.INIT_RAM_0C = 256'h060808082002102222800049323F1F003F0C0C31001C24102100202010000000;
defparam prom_inst_0.INIT_RAM_0D = 256'h02023F200000212104202012010208230200000000140220001404487F000800;
defparam prom_inst_0.INIT_RAM_0E = 256'h004104101004120C212221082021222121294920280408214020201120112155;
defparam prom_inst_0.INIT_RAM_0F = 256'h3E000400103F00214122427C3C2E00003C2E76104404185800103C3A3C5C3C00;
defparam prom_inst_0.INIT_RAM_10 = 256'h000408087F7F1022414962491248241E12121011241228103F1640401C611E19;
defparam prom_inst_0.INIT_RAM_11 = 256'h0C01004000001F1E083E3E220E04082504003F003F6302200008083E12000800;
defparam prom_inst_0.INIT_RAM_12 = 256'h0000040810080C0C212221081E3E223E212549203004083F403C3C11201E3F55;
defparam prom_inst_0.INIT_RAM_13 = 256'h3E000200200221124922421042311E3E42314910480008643E7C424642620200;
defparam prom_inst_0.INIT_RAM_14 = 256'h3008080820021022494914491208422112212012241230102129407824121125;
defparam prom_inst_0.INIT_RAM_15 = 256'h10023F20300001210821013F010808290800003000140220001510097F000800;
defparam prom_inst_0.INIT_RAM_16 = 256'h000004041010040C2D2221080128222021234120280408214720201120112156;
defparam prom_inst_0.INIT_RAM_17 = 256'h3E0004101004210C492242103020222142214910700408424210424240423E00;
defparam prom_inst_0.INIT_RAM_18 = 256'h49102A08100450144949083E1208422112211E14241228102109384024141F22;
defparam prom_inst_0.INIT_RAM_19 = 256'h1004001010300121082101020110083110000010002A02200022240912000000;
defparam prom_inst_0.INIT_RAM_1A = 256'h00000402102004122D22210801242A202123412024040821412020112011215C;
defparam prom_inst_0.INIT_RAM_1B = 256'h3E0004101008210C492242100C202221422149104804084242107E4240424200;
defparam prom_inst_0.INIT_RAM_1C = 256'h06201C0800003014494A14081208242212120118241225141209042024181125;
defparam prom_inst_0.INIT_RAM_1D = 256'h00080008100021210821210221200821200000100C49041000224A7E12000000;
defparam prom_inst_0.INIT_RAM_1E = 256'h0000040010200421331421082122262012214120224408212120201121112140;
defparam prom_inst_0.INIT_RAM_1F = 256'h3E00041010102312491442124220223142214910440408424610404642624600;
defparam prom_inst_0.INIT_RAM_20 = 256'h007E080800001036363C23080E08183C130C06103A33220C0C09181818101F19;
defparam prom_inst_0.INIT_RAM_21 = 256'h1810000420001E1E081E1E021E3F3E1E0018002000080808001D040812000800;
defparam prom_inst_0.INIT_RAM_22 = 256'h7F001C001C3F042121081E081E211D200C21413E21383E211E203F3E1E3E213E;
defparam prom_inst_0.INIT_RAM_23 = 256'h3E0038000E3F1D2136083C0C3C203E2E3C21490C42040C423A103E3A3C5C3B00;

endmodule //charROM
